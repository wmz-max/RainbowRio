`define TESTIO

`define UART_0_TX_DATA_ADDR 32'h0200_0000
`define UART_0_RX_DATA_ADDR 32'h0200_0001
`define UART_0_TX_CTRL_ADDR 32'h0200_0002
`define UART_0_TX_CTRL_ADDR 32'h0200_0003
`define UART_0_IRQ_PRIO_ADDR 32'h0200_0004
`define UART_0_IRQ_EN_ADDR 32'h0200_0005
`define UART_0_IRQ_IP_ADDR 32'h0200_0006
`define UART_1_TX_DATA_ADDR 32'h0200_0100
`define UART_1_RX_DATA_ADDR 32'h0200_0101
`define UART_1_TX_CTRL_ADDR 32'h0200_0102
`define UART_1_TX_CTRL_ADDR 32'h0200_0103
`define UART_1_IRQ_PRIO_ADDR 32'h0200_0104
`define UART_1_IRQ_EN_ADDR 32'h0200_0105
`define UART_1_IRQ_IP_ADDR 32'h0200_0106
`define UART_2_TX_DATA_ADDR 32'h0200_0200
`define UART_2_RX_DATA_ADDR 32'h0200_0201
`define UART_2_TX_CTRL_ADDR 32'h0200_0202
`define UART_2_TX_CTRL_ADDR 32'h0200_0203
`define UART_2_IRQ_PRIO_ADDR 32'h0200_0204
`define UART_2_IRQ_EN_ADDR 32'h0200_0205
`define UART_2_IRQ_IP_ADDR 32'h0200_0206
`define GPIO_SIZE 2
`define GPIO_0_VALUE_ADDR 32'h0200_0300
`define GPIO_0_INPUT_EN_ADDR 32'h0200_0301
`define GPIO_0_TX_OUTPUT_EN_ADDR 32'h0200_0302
`define GPIO_0_TX_PORT_ADDR 32'h0200_0303
`define GPIO_0_IRQ_PRIO_ADDR 32'h0200_0304
`define GPIO_0_IRQ_EN_ADDR 32'h0200_0305
`define GPIO_0_IRQ_IP_ADDR 32'h0200_0306
`define GPIO_1_VALUE_ADDR 32'h0200_0400
`define GPIO_1_INPUT_EN_ADDR 32'h0200_0401
`define GPIO_1_TX_OUTPUT_EN_ADDR 32'h0200_0402
`define GPIO_1_TX_PORT_ADDR 32'h0200_0403
`define GPIO_1_IRQ_PRIO_ADDR 32'h0200_0404
`define GPIO_1_IRQ_EN_ADDR 32'h0200_0405
`define GPIO_1_IRQ_IP_ADDR 32'h0200_0406
`define GPIO_2_VALUE_ADDR 32'h0200_0500
`define GPIO_2_INPUT_EN_ADDR 32'h0200_0501
`define GPIO_2_TX_OUTPUT_EN_ADDR 32'h0200_0502
`define GPIO_2_TX_PORT_ADDR 32'h0200_0503
`define GPIO_2_IRQ_PRIO_ADDR 32'h0200_0504
`define GPIO_2_IRQ_EN_ADDR 32'h0200_0505
`define GPIO_2_IRQ_IP_ADDR 32'h0200_0506
`define GPIO_3_VALUE_ADDR 32'h0200_0600
`define GPIO_3_INPUT_EN_ADDR 32'h0200_0601
`define GPIO_3_TX_OUTPUT_EN_ADDR 32'h0200_0602
`define GPIO_3_TX_PORT_ADDR 32'h0200_0603
`define GPIO_3_IRQ_PRIO_ADDR 32'h0200_0604
`define GPIO_3_IRQ_EN_ADDR 32'h0200_0605
`define GPIO_3_IRQ_IP_ADDR 32'h0200_0606
`define I2C_0_CMD_NOP_ADDR 32'h0200_0700
`define I2C_0_CMD_START_ADDR 32'h0200_0701
`define I2C_0_CMD_STOP_ADDR 32'h0200_0702
`define I2C_0_CMD_WRITE_ADDR 32'h0200_0703
`define I2C_0_CMD_READ_ADDR 32'h0200_0704
`define I2C_0_IRQ_PRIO_ADDR 32'h0200_0705
`define I2C_0_IRQ_EN_ADDR 32'h0200_0706
`define I2C_0_IRQ_IP_ADDR 32'h0200_0707
`define I2C_1_CMD_NOP_ADDR 32'h0200_0800
`define I2C_1_CMD_START_ADDR 32'h0200_0801
`define I2C_1_CMD_STOP_ADDR 32'h0200_0802
`define I2C_1_CMD_WRITE_ADDR 32'h0200_0803
`define I2C_1_CMD_READ_ADDR 32'h0200_0804
`define I2C_1_IRQ_PRIO_ADDR 32'h0200_0805
`define I2C_1_IRQ_EN_ADDR 32'h0200_0806
`define I2C_1_IRQ_IP_ADDR 32'h0200_0807
`define I2C_2_CMD_NOP_ADDR 32'h0200_0900
`define I2C_2_CMD_START_ADDR 32'h0200_0901
`define I2C_2_CMD_STOP_ADDR 32'h0200_0902
`define I2C_2_CMD_WRITE_ADDR 32'h0200_0903
`define I2C_2_CMD_READ_ADDR 32'h0200_0904
`define I2C_2_IRQ_PRIO_ADDR 32'h0200_0905
`define I2C_2_IRQ_EN_ADDR 32'h0200_0906
`define I2C_2_IRQ_IP_ADDR 32'h0200_0907
`define SPI_0_CFG_DATA_ADDR 32'h0200_0a00
`define SPI_0_IRQ_PRIO_ADDR 32'h0200_0a01
`define SPI_0_IRQ_EN_ADDR 32'h0200_0a02
`define SPI_0_IRQ_IP_ADDR 32'h0200_0a03
`define SPI_1_CFG_DATA_ADDR 32'h0200_0b00
`define SPI_1_IRQ_PRIO_ADDR 32'h0200_0b01
`define SPI_1_IRQ_EN_ADDR 32'h0200_0b02
`define SPI_1_IRQ_IP_ADDR 32'h0200_0b03
`define CORE_0_IRQ_TRSHD_ADDR 32'h0300_0000
`define CORE_0_IRQ_RESP_ADDR 32'h0300_0001
`define CORE_0_IRQ_COMP_ADDR 32'h0300_0002
`define CORE_1_IRQ_TRSHD_ADDR 32'h0300_0100
`define CORE_1_IRQ_RESP_ADDR 32'h0300_0101
`define CORE_1_IRQ_COMP_ADDR 32'h0300_0102
`define CORE_2_IRQ_TRSHD_ADDR 32'h0300_0200
`define CORE_2_IRQ_RESP_ADDR 32'h0300_0201
`define CORE_2_IRQ_COMP_ADDR 32'h0300_0202
`define CORE_3_IRQ_TRSHD_ADDR 32'h0300_0300
`define CORE_3_IRQ_RESP_ADDR 32'h0300_0301
`define CORE_3_IRQ_COMP_ADDR 32'h0300_0302
`define CORE_4_IRQ_TRSHD_ADDR 32'h0300_0400
`define CORE_4_IRQ_RESP_ADDR 32'h0300_0401
`define CORE_4_IRQ_COMP_ADDR 32'h0300_0402
localparam DEFAULT_FRENQUENCY = 50000000
localparam PERIPS_SIZE = 12
localparam WB_AD_WIDTH 43
localparam WB_DAT_WIDTH 32
localparam UART_CLK_FREQ 50000000
localparam CORE_NUM 5
localparam FREQUENCY1 = 50000000
localparam FREQUENCY2 = 50000000
localparam FREQUENCY3 = 50000000
localparam FREQUENCY4 = 50000000

